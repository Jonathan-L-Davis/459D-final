module top(
    input clk_100MHz_main, input isMealy_main, 
    input rst_main, input ctrl_input_main, 
    output reg clock_led,
    input [1:0] SW_input_main, 
    output [3:0] Anode_Activate_main,
    output [6:0] LED_out_main    
);


endmodule