module alucontrol(input [1:0] aluop, 
    input [5:0] funct, 
    output reg [2:0] alucont
    );

    always @(*) begin
        case(aluop)
            2'b00: alucont <= 3'b010; //add for lb/sb/addi
            2'b01: alucont <= 3'b110; //sub for beq
            default: case(funct)
                    6'b100000: alucont <= 3'b010; // add (for add)
                    6'b100010: alucont <= 3'b110; // subtract (for sub)
                    6'b100100: alucont <= 3'b000; // logical and (for and)
                    6'b100101: alucont <= 3'b001; // logical or (for or)
                    6'b101010: alucont <= 3'b111; // set on less (for slt)
                    default: alucont <= 3'b100; // should never happen
                endcase
        endcase
    end
endmodule
