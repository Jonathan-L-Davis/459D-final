module bus();
    // for part 3
endmodule